module %FILE% (
	%HERE%
);

%HERE%

endmodule

